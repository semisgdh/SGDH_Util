// timescale definition
`timescale 1ns/1ps